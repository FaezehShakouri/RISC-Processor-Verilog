`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:09:09 10/24/2020 
// Design Name: 
// Module Name:    Mux_16_to_1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: Using 4 to 1 mux and 2 to 1 mux.
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Mux_16_to_1();
	

endmodule
